/*###################################################################*\
##              Package Name:   param_pkg                            ##
##              Project Name: uart_tx_protocl                        ##
##              Date:   3/12/2023                                    ##
##              Author: Kholoud Ebrahim Darwseh                      ##
\*###################################################################*/

package param_pkg;
    parameter DWIDTH =6;
    parameter PERIOD = 5;
endpackage :param_pkg